// Engineer: Brett Duncan
//
// Create Date: 04/22/2023 05:06 PM


module alu_codes();

// // ALU Instructions
// localparam ADD = 3'h1;
// localparam SUB = 3'h2;
// localparam AND = 3'h3;
// localparam OR  = 3'h4;
// localparam SLL = 3'h5;
// localparam SRL = 3'h6;
// localparam NOP = 3'h0;

endmodule

