`include "alu.v"

module test_alu_subtract;

    initial begin
        $display("PASSED: test_alu_subtract");
    end

endmodule

